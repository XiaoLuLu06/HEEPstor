import TicSAT_pkg::*;

module TicSAT_FP32_Int8 #(
    parameter SA_SIZE = -1,

    // This parameters cannot be changed without recoding!!! They should be localparams,
    //  but DesignCompiler will complain. 

    parameter ACTIVATION_SIZE = 32
) (
    input logic resetn,
    input logic clk,

    // Used to load both weights and activations, depending on cmd
    input logic[ACTIVATION_SIZE-1:0] in_val,

    // Used to select in which FIFO position to write the input and read the output
    input logic[$clog2(SA_SIZE)-1:0] in_idx,

    output logic[ACTIVATION_SIZE-1:0] out,

    input command_t cmd
);

logic[ACTIVATION_SIZE-1:0] systolic_array_inputs[SA_SIZE-1:0];
logic[ACTIVATION_SIZE-1:0] systolic_array_outputs[SA_SIZE-1:0];

SA_FP32_Int8 #(
    .SA_SIZE            (SA_SIZE)
) u_SA_FP32_Int8 (
    .resetn             (resetn),
    .clk                (clk),
    .weight_input       (in_val),
    .inputs             (systolic_array_inputs),
    .outputs            (systolic_array_outputs),
    .cmd                (cmd)
);

FIFO_in #(
    .SA_SIZE            (SA_SIZE)
) u_FIFO_in (
    .resetn             (resetn),
    .clk                (clk),
    .in                 (in_val),
    .in_row_idx         (in_idx),
    .outputs            (systolic_array_inputs),
    .cmd                (cmd)
);

FIFO_out #(
    .SA_SIZE            (SA_SIZE)
) u_FIFO_out (
    .resetn             (resetn),
    .clk                (clk),
    .inputs             (systolic_array_outputs),
    .in_row_idx         (in_idx),
    .out                (out),
    .cmd                (cmd)
);

endmodule